`timescale 1ns / 1ps
/*
----------------------------------------------------------------------------------
--	(c) Rajesh Panicker
--	License terms :
--	You are free to use this code as long as you
--		(i) DO NOT post it on any public repository;
--		(ii) use it only for educational purposes;
--		(iii) accept the responsibility to ensure that your implementation does not violate any intellectual property of ARM Holdings or other entities.
--		(iv) accept that the program is provided "as is" without warranty of any kind or assurance regarding its suitability for any particular purpose;
--		(v) send an email to rajesh.panicker@ieee.org briefly mentioning its use (except when used for the course CG3207 at the National University of Singapore);
--		(vi) retain this notice in this file or any files derived from this.
----------------------------------------------------------------------------------
*/
module test_Wrapper #(
	   parameter N_LEDs_OUT	= 8,					
	   parameter N_DIPs		= 16,
	   parameter N_PBs		= 3 
	)
	(
	);
	
	// Signals for the Unit Under Test (UUT)
	reg  [N_DIPs-1:0] DIP = 0;		
	reg  [N_PBs-1:0] PB = 0;			
	wire [N_LEDs_OUT-1:0] LED_OUT;
	wire [6:0] LED_PC;			
	wire [31:0] SEVENSEGHEX;	
	wire [7:0] UART_TX;
	reg  UART_TX_ready = 0;
	wire UART_TX_valid;
	reg  [7:0] UART_RX = 0;
	reg  UART_RX_valid = 0;
	wire UART_RX_ack;
	wire OLED_Write;
	wire [6:0] OLED_Col;
	wire [5:0] OLED_Row;
	wire [23:0] OLED_Data;
	reg [31:0] ACCEL_Data;
	wire ACCEL_DReady;			
	reg  RESET = 0;	
	reg  CLK = 0;				
	
	// Instantiate UUT
    Wrapper dut(DIP, PB, LED_OUT, LED_PC, SEVENSEGHEX, UART_TX, UART_TX_ready, UART_TX_valid, UART_RX, UART_RX_valid, UART_RX_ack, OLED_Write, OLED_Col, OLED_Row, OLED_Data, ACCEL_Data, ACCEL_DReady, RESET, CLK) ;

	
	// Note: This testbench is for the Hello World program. Other assembly programs require appropriate modifications.
	// Run for about 6 us. Set UART_TX radix to ASCII to see the printed messages.
	// STIMULI
    initial
    begin
	RESET = 1; #10; RESET = 0; //hold reset state for 10 ns.
	    UART_TX_ready = 1'h1; // ok to keep it high continously in the testbench. In reality, it will be high only if UART is ready to send a data to PC
        UART_RX = 8'h50;// 'P'. Will be read and ignored by the processor
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack);
        wait(~UART_RX_ack);
        UART_RX_valid = 1'h0;
        #105;
        UART_RX = 8'h41;// 'A'
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack);
        wait(~UART_RX_ack);
	    UART_RX_valid = 1'h0;
        #105;
        UART_RX = 8'h0D;// '\r'
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack); // should print "Welcome to CG3207" following this.
        wait(~UART_RX_ack);
        UART_RX_valid = 1'h0;
        #2500
        // Run the simulation for about 3 us to see the full printed message. 
        
        // We are triggering a print one more time to see if it goes back correctly.
        // Run the simulation for another 3 us to see the full printed message a second time.
        
        UART_RX = 8'h50;// 'P'. Will be read and ignored by the processor
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack);
        wait(~UART_RX_ack);
        UART_RX_valid = 1'h0;
        #105;
        UART_RX = 8'h41;// 'A'
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack);
        wait(~UART_RX_ack);
	    UART_RX_valid = 1'h0;
        #105;
        UART_RX = 8'h0D;// '\r'
        UART_RX_valid = 1'h1;
        wait(UART_RX_ack); // should print "Welcome to CG3207" following this.
        wait(~UART_RX_ack);
        UART_RX_valid = 1'h0;
		//insert rest of the stimuli here
    end
	
	// GENERATE CLOCK       
    always          
    begin
       #5 CLK = ~CLK ; // invert clk every 5 time units 
    end
    
endmodule
